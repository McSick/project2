library ieee;
use ieee.std_logic_1164.all;
use ieee.NUMERIC_STD.all;
use ieee.std_logic_1164.STD_LOGIC;
entity mycpu is
		port ( 			
			CLK		:		in	std_logic;			
			nReset	:		in	std_logic;			
			halt	:		out	std_logic;
            ramAddr : out std_logic_vector(15 downto 0);
            ramData : out std_logic_vector(31 downto 0);
            ramWen  : out std_logic;
            ramRen  : out std_logic;
            ramQ    : in  std_logic_vector(31 downto 0);
            ramState : in std_logic_vector(1 downto 0)
		);	
	end mycpu;

architecture behavioral of mycpu is
  
   	component a32bitaddr 
  		port( A : in std_logic_vector(31 downto 0);
	      B : in std_logic_vector(31 downto 0);
	      SUM : out std_logic_vector(31 downto 0);
	      V : out std_logic);
	   end component;

	   component alu is
     port ( opcode:         IN STD_LOGIC_VECTOR (2 downto 0);
         A, B:           IN STD_LOGIC_VECTOR (31 downto 0);
         aluout:         OUT STD_LOGIC_VECTOR (31 downto 0);
         negative:       OUT STD_LOGIC;
         overflow, zero: OUT STD_LOGIC);
    end component;
      
	   component RegisterFile
	   port
	   (
		-- Write data input port
		wdat		:	in	std_logic_vector (31 downto 0);
		-- Select which register to write
		wsel		:	in	std_logic_vector (4 downto 0);
		-- Write Enable for entire register file
		wen			:	in	std_logic;
		-- clock, positive edge triggered
		clk			:	in	std_logic;
		-- REMEMBER: nReset-> '0' = RESET, '1' = RUN
		nReset	:	in	std_logic;
		-- Select which register to read on rdat1 
		rsel1		:	in	std_logic_vector (4 downto 0);
		-- Select which register to read on rdat2
		rsel2		:	in	std_logic_vector (4 downto 0);
		-- read port 1
		rdat1		:	out	std_logic_vector (31 downto 0);
		-- read port 2
		rdat2		:	out	std_logic_vector (31 downto 0)
		);
		end component;

		component  Extender
		 port(
    Instruction : in std_logic_vector(15 downto 0);
    ExtType : in std_logic;
    Im32 : out std_logic_vector(31 downto 0));
end component;
  	    
 	component SSC is
  port(
    opcode : in std_logic_vector(5 downto 0);
    funct : in std_logic_vector(5 downto 0);
    ExtType : out std_logic;
    WriteEnable : out std_logic;
    RegDst : out std_logic;
    AluSrc : out std_logic;
    ALU_cntrl : out std_logic_vector(2 downto 0);
    MemWrite : out std_logic; 
    MemOut : out std_logic;
    Branch : out std_logic;
    Jump : out std_logic;
    BNE : out std_logic;
    LUI :out std_logic

  );
end component;


component pipeline_controller IS
	PORT
	(
		memstate	: IN STD_LOGIC;
		ExC			: OUT STD_LOGIC;
		WBC			: OUT STD_LOGIC;
		MEMC		: OUT STD_LOGIC;	
		IDC			: OUT STD_LOGIC
	);
end component;

  signal PC,Instruction,MemoryData : std_logic_vector(31 downto 0);

--Internal Signal declarations
signal memoryAddress : std_logic_vector(15 downto 0);

signal ExtType,memwait,nResetSynch : std_logic;
signal WriteEnable : std_logic;
signal RegDst : std_logic;
signal AluSrc : std_logic;
signal ALUcntr : std_logic_vector(2 downto 0);
signal MemWrite,MemOutMux,lui : std_logic;
signal Branch : std_logic;
signal Jump,HaltI,BNE : std_logic;
Signal WriteDataReg : std_logic_vector(31 downto 0);
signal zero,overflow,over1,over2 : std_logic;
signal negative : std_logic;
signal BusA, BusB,Im32,Bsel,PCP4,PCJmp,PCJmp_stg4,JumpAddress,BranchAddress,AlmostPCnextPC,ALUout,shifted,WriteDataReg2: std_logic_vector(31 downto 0);
signal rs,rt,rd,rtd : std_logic_vector(4 downto 0);
signal memstate : std_logic;
-- Stage 1
-- Stage 2
signal PCP4_stg2, Instruction_stg2 : std_logic_vector(31 downto 0);
signal memstate_stg2,Stall_23 : std_logic;
signal ExC,WBC,MEMC :std_logic;
-- Stage 3
signal BusA_stg3,BusB_stg3,PCP4_stg3, Instruction_stg3 : std_logic_vector(31 downto 0);
signal ExC_stg3,WBC_stg3,MEMC_stg3 :std_logic;
-- Stage 4
signal Instruction_stg4 : std_logic_vector(31 downto 0);
signal zero_stg4
-- Stage 5
signal Instruction_stg5 : std_logic_vector(31 downto 0);

TYPE STATE_TYPE IS (s0 ,s1);
  Signal state,nextstate : STATE_TYPE;

begin

		imemAddr <= PC;
		imemData <= Instruction;
		dmemDataRead <= MemoryData;
		dmemDataWrite <= BusB;
         
    dmemAddr <= ALUout;
  
  rd <= Instruction_stg3(15 downto 11);
  rt <= Instruction_stg3(20 downto 16);
  rs <= Instruction(25 downto 21);
  
  --Mux Regdst
  with RegDst select
    rtd <= rd when '1', rt when '0',"00000" when others;
    
    
  ExBlock : Extender
  Port map(Instruction_stg2(15 downto 0),ExtType,Im32);
  
  
  --Mux AluSrc
  with AluSrc select
    BSel <= Im32_stg3 when '1', BusB_stg3 when others;
    
   AluBlock : alu
   Port map(ALUcntr,BusA_stg3,Bsel,ALUout,negative, overflow,zero);
 

   
   
   with MemOutMux select
    WriteDataReg <= ALUout when '1', MemoryData when others;
    
    
    with lui select
    WriteDataReg2 <= Instruction(15 downto 0) & x"0000" when  '1', WriteDataReg when others;
    
    
  RegisterBlock : registerFile
  Port map(WriteDataReg2,rtd,WriteEnable,clk,nReset,rs,rt,BusA,BusB);
  
  ControllerBlock : SSC
  Port map(Instruction(31 downto 26),Instruction(5 downto 0),ExtType,WriteEnable,RegDst,AluSrc,ALUcntr,MemWrite,MemOutMux,Branch,Jump,BNE,lui);
 
branchand :  process(Instruction)
begin
  IF(Instruction_stg5 = x"FFFFFFFF") then
  HaltI <= '1';
else
  HaltI <= '0';
end if;
end process;
  
  
twocycle : process(clk,nReset)
begin
  if(nReset = '0') then
    state <= s0;
elsif(rising_edge(CLK)) then
  state <= nextstate;
end if;
end process;

twocycleo : process(state,Instruction)
begin
  case state is
  when s0 =>
     IF(Instruction(31 downto 26) = "100011") then
    nextstate <= s1;
    memwait <= '1';
  else
    memwait <= '0';
    nextstate <= s0;
  end if;
   when s1 =>
   nextstate <= s0;
   memwait <= '0';
   end case;
end process;
 
 Halt <= HaltI;
 with (HaltI or memwait) select
    NextPC <= PC when '1', AlmostPC when others;
    
  
  ADDPC4 : a32bitaddr
  Port map(PC,x"00000004",PCP4,over1);
    
  shifted <=Im32_stg3(29 downto 0) & "00";
    
  ADDBR : a32bitaddr
  Port map(PCP4_stg3,shifted, PCJmp,over2);
    
  
  with ((Branch AND zero_stg4) or (BNE AND (not zero_stg4))) select
   BranchAddress <= PCJmp_stg4 when '1', PCP4_stg4 when others;
   
   with Jump select
    AlmostPC <= PCP4_stg4(31 downto 28) & Instruction_stg4(25 downto 0) & "00" when '1', BranchAddress when others;
    
     registers : process (CLK, nReset,nResetSynch)
     begin
         if (nReset = '0') then		 
		-- Reset here		
		PC <= x"00000000";
	 elsif (rising_edge(CLK))and(Stall = '0') then
		if(nResetSynch = '0') then
			PC <= x"00000000";
		else		
			PC <= nextPC;
		end if;
	end if;       
     end process;
     IFIDRegister: process(CLK,nReset,nResetSynch_S12,Stall_S45)		--Stage 1-2
	begin
	if (nReset = '0') then
		memstate_stg2 <= '0';
		Instruction_stg2 <=  x"00000000";
		PCP4_stg2 <= x"00000000";
	elsif (rising_edge(CLK))and(Stall = '0') then
		if(nResetSynch = '0') then
			memstate_stg2 <= '0';
			Instruction_stg2 <=  x"00000000";
			PCP4_stg2 <= x"00000000";
		else
			memstate_stg2 <= memstate;
			Instruction_stg2 <= Instruction;
			PCP4_stg2 <= PCP4;				
		end if;
	end if;
     end process;
     IDEXRegister: process(CLK,nReset,nResetSynch_S23,Stall_S45)		--Stage 2-3
	begin
	if (nReset = '0') then
		BusA_stg3 <= "00000";
	 	BusB_stg3 <= "00000";
		Im32_stg3 <= x"00000000";
		ExC_stg3 <= x"00";
		WBC_stg3 <= x"00";				
		MEMC_stg3 <= x"00";		
		Instruction_stg3 <=  x"00000000";		
		PCP4_stg3 <=  x"00000000";
	elsif (rising_edge(CLK))and(Stall = '0') then
		if(nResetSynch = '0') then
			BusA_stg3 <= "00000";
		 	BusB_stg3 <= "00000";
			Im32_stg3 <= x"00000000";
			ExC_stg3 <= x"00";
			WBC_stg3 <= x"00";				
			MEMC_stg3 <= x"00";		
			Instruction_stg3 <=  x"00000000";		
			PCP4_stg3 <=  x"00000000";
		else
			BusA_stg3 <= BusA;
		 	BusB_stg3 <= BusB;
			Im32_stg3 <= Im32;
			ExC_stg3 <= ExC;
			WBC_stg3 <= WBC;
			MEMC_stg3 <= MEMC;
			Instruction_stg3 <= Instruction_stg2;
			PCP4_stg3 <= PCP4_stg2;
		end if;
	end if;
     end process;
     EXMEMRegister: process(CLK,nReset,nResetSynch_S34,Stall_S45)		--Stage 3-4
	begin
	if (nReset = '0') then
		PCP4_stg4 <= x"00000000";
		zero_stg4 <= '0';
		WBC_stg4 <= "00";
		Instruction_stg4 <=  x"00000000";
		MEMC_stg4 <= x"000";
	elsif (rising_edge(CLK))and(Stall = '0') then
		if(nResetSynch = '0') then
			PCP4_stg4 <= x"00000000";
			zero_stg4 <= '0';
			WBC_stg4 <= "00";
			Instruction_stg4 <=  x"00000000";
			MEMC_stg4 <= x"000";
		else
			PCP4_stg4 <= PCP4_stg3;
			zero_stg4 <= zero;
			WBC_stg4 <= WBC_stg3;
			Instruction_stg4 <= Instruction_stg3;
			MEMC_stg4 <= MEM3;
		end if;
	end if;
     end process;
     MEMWBRegister: process(CLK,nReset,nResetSynch_S45,Stall_S45)		--Stage 4-5
	begin
	if (nReset = '0') then
		WBC_stg5 <= WBC_stg4;
		Instruction_stg5 <=  x"00000000";
	elsif (rising_edge(CLK))and(Stall = '0') then
		if(nResetSynch = '0') then
			WBC_stg5 <= WBC_stg4;
			Instruction_stg5 <=  x"00000000";
		else
			WBC_stg5 <= WBC_stg4;															
			Instruction_stg5 <= Instruction_stg4;
		end if;
	end if;
     end process;
     
     with haltI select
      memoryAddress <= dumpAddr when '1',ALUout(15 downto 0) when others;
      

      
 
    --RAM D
  DataMemory : ramd
	PORT Map	(memoryAddress,CLK,BusB,MemWrite,MemoryData);

  InstructionMemory : rami
  Port map (PC(15 downto 0),CLK,PC,'0',Instruction);
  
  PipelineController: pipeline_controller
	PORT Map (memstate_stg2,ExC,WBC,MEMC,IDC);
  

  
end behavioral;
